library ieee;
use ieee.std_logic_1164.all;

entity EN_MUX41_cond is 
  port (
    A, B, C, D : in  std_logic;
    S0, S1     : in  std_logic;
    Y          : out std_logic
  );
end EN_MUX41_cond;

architecture RTL of EN_MUX41_cond is
begin
  -- S1 S0: 00->A, 01->B, 10->C, 11->D
  Y <= A when (S1 = '0' and S0 = '0') else
       B when (S1 = '0' and S0 = '1') else
       C when (S1 = '1' and S0 = '0') else
       D when (S1 = '1' and S0 = '1') else
       'X'; -- fallback for non '0'/'1' on selects
end RTL;